ֻ���Ƿ�֧b,����������˷�֧�b�Ĺ����
