����һ���µ��ļ����з�֧a�����������˷�֧a���¹���
